`include "driver.sv"
`include "environment.sv"
`include "monitor.sv"
`include "tb_top.sv"
`include "ahp.v"
`include "ahp_tb.v"
